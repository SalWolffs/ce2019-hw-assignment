-- unclocked ROM containing VLIW instructions from page 9
-- generated with python

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity rbc_rom is
    generic(
        ws: integer := 18;
        ads: integer := 7);
    port(
        address: in std_logic_vector(ads-1 downto 0);
        dout: out std_logic_vector(ws-1 downto 0));
end rbc_rom;

architecture behavioral of rbc_rom is
type rom is array(0 to 2**ads-1) of std_logic_vector(ws-1 downto 0);
constant data: rom := (
    000 => "001011000001100110",
    001 => "001011010010000111",
    002 => "001011100010101000",
    003 => "010011110001100100",
    004 => "010100000011000111",
    005 => "001011110111110000",
    006 => "010100000110001101",
    007 => "011011110111110000",
    008 => "010100000010000101",
    009 => "010100010011101000",
    010 => "001100001000010001",
    011 => "010100010110101110",
    012 => "011100001000010001",
    013 => "010100010001100101",
    014 => "010100100011001000",
    015 => "001100011000110010",
    016 => "010100100110001110",
    017 => "011100101000110010",
    018 => "001100110001001110",
    019 => "011100011001010011",
    020 => "010100111000110001",
    021 => "010100011000110011",
    022 => "011100110110110001",
    023 => "010100010110110001",
    024 => "001100100001010010",
    025 => "010011010111001110",
    026 => "010011100110101110",
    027 => "011100101001001110",
    028 => "011100101001001100",
    029 => "010011011001010010",
    030 => "010100100110110010",
    031 => "010011010110001100",
    032 => "010011000110101100",
    033 => "011011000110001110",
    034 => "001011011000010010",
    035 => "001011100110010010",
    036 => "001100101000110011",
    037 => "010010101001001110",
    038 => "001100010111110001",
    039 => "011010011000101101",
    040 => "001100111000010011",
    041 => "001011010111101100",
    042 => "010010111001101101",
    043 => "000000000000000000",
    044 => "001011000001100011",
    045 => "001011010010000100",
    046 => "001011100010100101",
    047 => "001011110001100100",
    048 => "010011110111101111",
    049 => "001100100001100101",
    050 => "010100101001010010",
    051 => "001100010001001110",
    052 => "011100011000110010",
    053 => "010100001000110001",
    054 => "010100011000010001",
    055 => "011100000110110001",
    056 => "010100010110110001",
    057 => "001100011000010001",
    058 => "001100001000001111",
    059 => "010011110111001110",
    060 => "010011100111001111",
    061 => "001100100001010010",
    062 => "011100101001001110",
    063 => "011100101001001100",
    064 => "010011111001010010",
    065 => "010100101001001111",
    066 => "010011110110001100",
    067 => "010011000111101100",
    068 => "011011000110001110",
    069 => "001011000110010010",
    070 => "001011100010000101",
    071 => "010011100111001110",
    072 => "010010101000101100",
    073 => "001100100111010010",
    074 => "011010011000010010",
    075 => "001100100111001101",
    076 => "010100101001010010",
    077 => "010010111001010010",
    078 => "000000000000000000",
    079 => "000000000000000000",
    080 => "000000000000000000",
    081 => "000000000000000000",
    082 => "000000000000000000",
    083 => "000000000000000000",
    084 => "000000000000000000",
    085 => "000000000000000000",
    086 => "000000000000000000",
    087 => "000000000000000000",
    088 => "000000000000000000",
    089 => "000000000000000000",
    090 => "000000000000000000",
    091 => "000000000000000000",
    092 => "000000000000000000",
    093 => "000000000000000000",
    094 => "000000000000000000",
    095 => "000000000000000000",
    096 => "000000000000000000",
    097 => "000000000000000000",
    098 => "000000000000000000",
    099 => "000000000000000000",
    100 => "000000000000000000",
    101 => "000000000000000000",
    102 => "000000000000000000",
    103 => "000000000000000000",
    104 => "000000000000000000",
    105 => "000000000000000000",
    106 => "000000000000000000",
    107 => "000000000000000000",
    108 => "000000000000000000",
    109 => "000000000000000000",
    110 => "000000000000000000",
    111 => "000000000000000000",
    112 => "000000000000000000",
    113 => "000000000000000000",
    114 => "000000000000000000",
    115 => "000000000000000000",
    116 => "000000000000000000",
    117 => "000000000000000000",
    118 => "000000000000000000",
    119 => "000000000000000000",
    120 => "000000000000000000",
    121 => "000000000000000000",
    122 => "000000000000000000",
    123 => "000000000000000000",
    124 => "000000000000000000",
    125 => "000000000000000000",
    126 => "000000000000000000",
    127 => "000000000000000000");

begin
    dout <= data(to_integer(to_01(unsigned(address))));
end behavioral;
