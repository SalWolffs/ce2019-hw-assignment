-- unclocked ROM containing VLIW instructions from page 9
-- generated with python

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity rbc_rom is
    generic(
        ws: integer := 18;
        ads: integer := 7);
    port(
        address: in std_logic_vector(ads-1 downto 0);
        dout: out std_logic_vector(ws-1 downto 0));
end rbc_rom;

architecture behavioral of rbc_rom is
type rom is array(0 to 2**ads-1) of std_logic_vector(ws-1 downto 0);
constant data: rom := (
    000 => "100000000000000000",
    001 => "001011000011000011",
    002 => "001011010011100100",
    003 => "001011100100000101",
    004 => "010011110010000011",
    005 => "010100000011100110",
    006 => "001011111000001111",
    007 => "010100000110101100",
    008 => "011011111000001111",
    009 => "010100000010100100",
    010 => "010100010100000111",
    011 => "001100001000110000",
    012 => "010100010111001101",
    013 => "011100001000110000",
    014 => "010100010010100011",
    015 => "010100100100000110",
    016 => "001100011001010001",
    017 => "010100100111001100",
    018 => "011100101001010001",
    019 => "001100110111000010",
    020 => "011100011001110010",
    021 => "010100111000110001",
    022 => "010100011001110001",
    023 => "011100111000101101",
    024 => "010100011000101101",
    025 => "001100101001000010",
    026 => "010011010111001110",
    027 => "010011100111001101",
    028 => "011100100111010010",
    029 => "011100100110010010",
    030 => "010011011001010010",
    031 => "010100101001001101",
    032 => "010011010110001100",
    033 => "010011000110001101",
    034 => "011011000111001100",
    035 => "001011011001010000",
    036 => "001011101001001100",
    037 => "001100101001110001",
    038 => "010010100111010010",
    039 => "001100011000101111",
    040 => "011010010110110001",
    041 => "001100111001110000",
    042 => "001011010110001111",
    043 => "010010110110110011",
    044 => "000000000000000000",
    045 => "100000000000000000",
    046 => "001011000001100011",
    047 => "001011010010000100",
    048 => "001011100010100101",
    049 => "001011110010000011",
    050 => "010011110111101111",
    051 => "001100100010100011",
    052 => "010100101001010010",
    053 => "001100010111000010",
    054 => "011100011001010001",
    055 => "010100001000110001",
    056 => "010100011000110000",
    057 => "011100001000101101",
    058 => "010100011000101101",
    059 => "001100011000110000",
    060 => "001100000111110000",
    061 => "010011110111001110",
    062 => "010011100111101110",
    063 => "001100101001000010",
    064 => "011100100111010010",
    065 => "011100100110010010",
    066 => "010011111001010010",
    067 => "010100100111110010",
    068 => "010011110110001100",
    069 => "010011000110001111",
    070 => "011011000111001100",
    071 => "001011001001001100",
    072 => "001011100010100100",
    073 => "010011100111001110",
    074 => "010010100110010001",
    075 => "001100101001001110",
    076 => "011010011001010000",
    077 => "001100100110101110",
    078 => "010100101001010010",
    079 => "010010111001010010",
    080 => "000000000000000000",
    081 => "000000000000000000",
    082 => "000000000000000000",
    083 => "000000000000000000",
    084 => "000000000000000000",
    085 => "000000000000000000",
    086 => "000000000000000000",
    087 => "000000000000000000",
    088 => "000000000000000000",
    089 => "000000000000000000",
    090 => "000000000000000000",
    091 => "000000000000000000",
    092 => "000000000000000000",
    093 => "000000000000000000",
    094 => "000000000000000000",
    095 => "000000000000000000",
    096 => "000000000000000000",
    097 => "000000000000000000",
    098 => "000000000000000000",
    099 => "000000000000000000",
    100 => "000000000000000000",
    101 => "000000000000000000",
    102 => "000000000000000000",
    103 => "000000000000000000",
    104 => "000000000000000000",
    105 => "000000000000000000",
    106 => "000000000000000000",
    107 => "000000000000000000",
    108 => "000000000000000000",
    109 => "000000000000000000",
    110 => "000000000000000000",
    111 => "000000000000000000",
    112 => "000000000000000000",
    113 => "000000000000000000",
    114 => "000000000000000000",
    115 => "000000000000000000",
    116 => "000000000000000000",
    117 => "000000000000000000",
    118 => "000000000000000000",
    119 => "000000000000000000",
    120 => "000000000000000000",
    121 => "000000000000000000",
    122 => "000000000000000000",
    123 => "000000000000000000",
    124 => "000000000000000000",
    125 => "000000000000000000",
    126 => "000000000000000000",
    127 => "000000000000000000");

begin
    dout <= data(to_integer(to_01(unsigned(address))));
end behavioral;
